module regfile(
    input logic clock,
    input logic [4:0] read_address_0,
    input logic [4:0] read_address_1,
    input logic [4:0] write_address_0,
    input logic write_enable_0,
    input logic [31:0] write_data_0,
    output logic [31:0] read_data_0,
    output logic [31:0] read_data_1
);

logic [31:0] conditionalnode$0;
assign read_data_0 = conditionalnode$0;

logic [31:0] conditionalnode$1;
assign read_data_1 = conditionalnode$1;

logic eqnode$2;
logic [31:0] repeatnode$3;
logic [31:0] conditionalnode$4;
assign conditionalnode$0 = eqnode$2 ? repeatnode$3 : conditionalnode$4;

logic eqnode$5;
logic [31:0] repeatnode$6;
logic [31:0] conditionalnode$7;
assign conditionalnode$1 = eqnode$5 ? repeatnode$6 : conditionalnode$7;

logic [4:0] wirenode$8;
logic [4:0] zeroextendnode$9;
assign eqnode$2 = wirenode$8 == zeroextendnode$9;

assign repeatnode$3 = {32{1'b0}};

logic andnode$10;
logic [31:0] wirenode$11;
logic [31:0] conditionalnode$12;
assign conditionalnode$4 = andnode$10 ? wirenode$11 : conditionalnode$12;

logic [4:0] wirenode$13;
logic [4:0] zeroextendnode$14;
assign eqnode$5 = wirenode$13 == zeroextendnode$14;

assign repeatnode$6 = {32{1'b0}};

logic andnode$15;
logic [31:0] conditionalnode$16;
assign conditionalnode$7 = andnode$15 ? wirenode$11 : conditionalnode$16;

assign wirenode$8 = read_address_0;

assign zeroextendnode$9 = '0;

logic eqnode$17;
logic wirenode$18;
assign andnode$10 = eqnode$17 & wirenode$18;

assign wirenode$11 = write_data_0;

logic eqnode$19;
logic [31:0] registernode$20;
logic [31:0] conditionalnode$21;
assign conditionalnode$12 = eqnode$19 ? registernode$20 : conditionalnode$21;

assign wirenode$13 = read_address_1;

assign zeroextendnode$14 = '0;

logic eqnode$22;
assign andnode$15 = eqnode$22 & wirenode$18;

logic eqnode$23;
logic [31:0] conditionalnode$24;
assign conditionalnode$16 = eqnode$23 ? registernode$20 : conditionalnode$24;

logic [4:0] wirenode$25;
assign eqnode$17 = wirenode$8 == wirenode$25;

assign wirenode$18 = write_enable_0;

logic [4:0] zeroextendnode$26;
assign eqnode$19 = wirenode$8 == zeroextendnode$26;

logic [31:0] wirenode$27;
always_ff @ (posedge clock) registernode$20 <= wirenode$27;

logic eqnode$28;
logic [31:0] registernode$29;
logic [31:0] conditionalnode$30;
assign conditionalnode$21 = eqnode$28 ? registernode$29 : conditionalnode$30;

assign eqnode$22 = wirenode$13 == wirenode$25;

logic [4:0] zeroextendnode$31;
assign eqnode$23 = wirenode$13 == zeroextendnode$31;

logic eqnode$32;
logic [31:0] conditionalnode$33;
assign conditionalnode$24 = eqnode$32 ? registernode$29 : conditionalnode$33;

assign wirenode$25 = write_address_0;

assign zeroextendnode$26 = 1'b1;

logic [31:0] conditionalnode$34;
assign wirenode$27 = conditionalnode$34;

logic [4:0] zeroextendnode$35;
assign eqnode$28 = wirenode$8 == zeroextendnode$35;

logic [31:0] wirenode$36;
always_ff @ (posedge clock) registernode$29 <= wirenode$36;

logic eqnode$37;
logic [31:0] registernode$38;
logic [31:0] conditionalnode$39;
assign conditionalnode$30 = eqnode$37 ? registernode$38 : conditionalnode$39;

assign zeroextendnode$31 = 1'b1;

logic [4:0] zeroextendnode$40;
assign eqnode$32 = wirenode$13 == zeroextendnode$40;

logic eqnode$41;
logic [31:0] conditionalnode$42;
assign conditionalnode$33 = eqnode$41 ? registernode$38 : conditionalnode$42;

logic andnode$43;
assign conditionalnode$34 = andnode$43 ? wirenode$11 : registernode$20;

assign zeroextendnode$35 = 2'b10;

logic [31:0] conditionalnode$44;
assign wirenode$36 = conditionalnode$44;

logic [4:0] zeroextendnode$45;
assign eqnode$37 = wirenode$8 == zeroextendnode$45;

logic [31:0] wirenode$46;
always_ff @ (posedge clock) registernode$38 <= wirenode$46;

logic eqnode$47;
logic [31:0] registernode$48;
logic [31:0] conditionalnode$49;
assign conditionalnode$39 = eqnode$47 ? registernode$48 : conditionalnode$49;

assign zeroextendnode$40 = 2'b10;

logic [4:0] zeroextendnode$50;
assign eqnode$41 = wirenode$13 == zeroextendnode$50;

logic eqnode$51;
logic [31:0] conditionalnode$52;
assign conditionalnode$42 = eqnode$51 ? registernode$48 : conditionalnode$52;

logic eqnode$53;
assign andnode$43 = eqnode$53 & wirenode$18;

logic andnode$54;
assign conditionalnode$44 = andnode$54 ? wirenode$11 : registernode$29;

assign zeroextendnode$45 = 2'b11;

logic [31:0] conditionalnode$55;
assign wirenode$46 = conditionalnode$55;

logic [4:0] zeroextendnode$56;
assign eqnode$47 = wirenode$8 == zeroextendnode$56;

logic [31:0] wirenode$57;
always_ff @ (posedge clock) registernode$48 <= wirenode$57;

logic eqnode$58;
logic [31:0] registernode$59;
logic [31:0] conditionalnode$60;
assign conditionalnode$49 = eqnode$58 ? registernode$59 : conditionalnode$60;

assign zeroextendnode$50 = 2'b11;

logic [4:0] zeroextendnode$61;
assign eqnode$51 = wirenode$13 == zeroextendnode$61;

logic eqnode$62;
logic [31:0] conditionalnode$63;
assign conditionalnode$52 = eqnode$62 ? registernode$59 : conditionalnode$63;

logic [4:0] zeroextendnode$64;
assign eqnode$53 = wirenode$25 == zeroextendnode$64;

logic eqnode$65;
assign andnode$54 = eqnode$65 & wirenode$18;

logic andnode$66;
assign conditionalnode$55 = andnode$66 ? wirenode$11 : registernode$38;

assign zeroextendnode$56 = 3'b100;

logic [31:0] conditionalnode$67;
assign wirenode$57 = conditionalnode$67;

logic [4:0] zeroextendnode$68;
assign eqnode$58 = wirenode$8 == zeroextendnode$68;

logic [31:0] wirenode$69;
always_ff @ (posedge clock) registernode$59 <= wirenode$69;

logic eqnode$70;
logic [31:0] registernode$71;
logic [31:0] conditionalnode$72;
assign conditionalnode$60 = eqnode$70 ? registernode$71 : conditionalnode$72;

assign zeroextendnode$61 = 3'b100;

logic [4:0] zeroextendnode$73;
assign eqnode$62 = wirenode$13 == zeroextendnode$73;

logic eqnode$74;
logic [31:0] conditionalnode$75;
assign conditionalnode$63 = eqnode$74 ? registernode$71 : conditionalnode$75;

assign zeroextendnode$64 = 1'b1;

logic [4:0] zeroextendnode$76;
assign eqnode$65 = wirenode$25 == zeroextendnode$76;

logic eqnode$77;
assign andnode$66 = eqnode$77 & wirenode$18;

logic andnode$78;
assign conditionalnode$67 = andnode$78 ? wirenode$11 : registernode$48;

assign zeroextendnode$68 = 3'b101;

logic [31:0] conditionalnode$79;
assign wirenode$69 = conditionalnode$79;

logic [4:0] zeroextendnode$80;
assign eqnode$70 = wirenode$8 == zeroextendnode$80;

logic [31:0] wirenode$81;
always_ff @ (posedge clock) registernode$71 <= wirenode$81;

logic eqnode$82;
logic [31:0] registernode$83;
logic [31:0] conditionalnode$84;
assign conditionalnode$72 = eqnode$82 ? registernode$83 : conditionalnode$84;

assign zeroextendnode$73 = 3'b101;

logic [4:0] zeroextendnode$85;
assign eqnode$74 = wirenode$13 == zeroextendnode$85;

logic eqnode$86;
logic [31:0] conditionalnode$87;
assign conditionalnode$75 = eqnode$86 ? registernode$83 : conditionalnode$87;

assign zeroextendnode$76 = 2'b10;

logic [4:0] zeroextendnode$88;
assign eqnode$77 = wirenode$25 == zeroextendnode$88;

logic eqnode$89;
assign andnode$78 = eqnode$89 & wirenode$18;

logic andnode$90;
assign conditionalnode$79 = andnode$90 ? wirenode$11 : registernode$59;

assign zeroextendnode$80 = 3'b110;

logic [31:0] conditionalnode$91;
assign wirenode$81 = conditionalnode$91;

logic [4:0] zeroextendnode$92;
assign eqnode$82 = wirenode$8 == zeroextendnode$92;

logic [31:0] wirenode$93;
always_ff @ (posedge clock) registernode$83 <= wirenode$93;

logic eqnode$94;
logic [31:0] registernode$95;
logic [31:0] conditionalnode$96;
assign conditionalnode$84 = eqnode$94 ? registernode$95 : conditionalnode$96;

assign zeroextendnode$85 = 3'b110;

logic [4:0] zeroextendnode$97;
assign eqnode$86 = wirenode$13 == zeroextendnode$97;

logic eqnode$98;
logic [31:0] conditionalnode$99;
assign conditionalnode$87 = eqnode$98 ? registernode$95 : conditionalnode$99;

assign zeroextendnode$88 = 2'b11;

logic [4:0] zeroextendnode$100;
assign eqnode$89 = wirenode$25 == zeroextendnode$100;

logic eqnode$101;
assign andnode$90 = eqnode$101 & wirenode$18;

logic andnode$102;
assign conditionalnode$91 = andnode$102 ? wirenode$11 : registernode$71;

assign zeroextendnode$92 = 3'b111;

logic [31:0] conditionalnode$103;
assign wirenode$93 = conditionalnode$103;

logic [4:0] zeroextendnode$104;
assign eqnode$94 = wirenode$8 == zeroextendnode$104;

logic [31:0] wirenode$105;
always_ff @ (posedge clock) registernode$95 <= wirenode$105;

logic eqnode$106;
logic [31:0] registernode$107;
logic [31:0] conditionalnode$108;
assign conditionalnode$96 = eqnode$106 ? registernode$107 : conditionalnode$108;

assign zeroextendnode$97 = 3'b111;

logic [4:0] zeroextendnode$109;
assign eqnode$98 = wirenode$13 == zeroextendnode$109;

logic eqnode$110;
logic [31:0] conditionalnode$111;
assign conditionalnode$99 = eqnode$110 ? registernode$107 : conditionalnode$111;

assign zeroextendnode$100 = 3'b100;

logic [4:0] zeroextendnode$112;
assign eqnode$101 = wirenode$25 == zeroextendnode$112;

logic eqnode$113;
assign andnode$102 = eqnode$113 & wirenode$18;

logic andnode$114;
assign conditionalnode$103 = andnode$114 ? wirenode$11 : registernode$83;

assign zeroextendnode$104 = 4'b1000;

logic [31:0] conditionalnode$115;
assign wirenode$105 = conditionalnode$115;

logic [4:0] zeroextendnode$116;
assign eqnode$106 = wirenode$8 == zeroextendnode$116;

logic [31:0] wirenode$117;
always_ff @ (posedge clock) registernode$107 <= wirenode$117;

logic eqnode$118;
logic [31:0] registernode$119;
logic [31:0] conditionalnode$120;
assign conditionalnode$108 = eqnode$118 ? registernode$119 : conditionalnode$120;

assign zeroextendnode$109 = 4'b1000;

logic [4:0] zeroextendnode$121;
assign eqnode$110 = wirenode$13 == zeroextendnode$121;

logic eqnode$122;
logic [31:0] conditionalnode$123;
assign conditionalnode$111 = eqnode$122 ? registernode$119 : conditionalnode$123;

assign zeroextendnode$112 = 3'b101;

logic [4:0] zeroextendnode$124;
assign eqnode$113 = wirenode$25 == zeroextendnode$124;

logic eqnode$125;
assign andnode$114 = eqnode$125 & wirenode$18;

logic andnode$126;
assign conditionalnode$115 = andnode$126 ? wirenode$11 : registernode$95;

assign zeroextendnode$116 = 4'b1001;

logic [31:0] conditionalnode$127;
assign wirenode$117 = conditionalnode$127;

logic [4:0] zeroextendnode$128;
assign eqnode$118 = wirenode$8 == zeroextendnode$128;

logic [31:0] wirenode$129;
always_ff @ (posedge clock) registernode$119 <= wirenode$129;

logic eqnode$130;
logic [31:0] registernode$131;
logic [31:0] conditionalnode$132;
assign conditionalnode$120 = eqnode$130 ? registernode$131 : conditionalnode$132;

assign zeroextendnode$121 = 4'b1001;

logic [4:0] zeroextendnode$133;
assign eqnode$122 = wirenode$13 == zeroextendnode$133;

logic eqnode$134;
logic [31:0] conditionalnode$135;
assign conditionalnode$123 = eqnode$134 ? registernode$131 : conditionalnode$135;

assign zeroextendnode$124 = 3'b110;

logic [4:0] zeroextendnode$136;
assign eqnode$125 = wirenode$25 == zeroextendnode$136;

logic eqnode$137;
assign andnode$126 = eqnode$137 & wirenode$18;

logic andnode$138;
assign conditionalnode$127 = andnode$138 ? wirenode$11 : registernode$107;

assign zeroextendnode$128 = 4'b1010;

logic [31:0] conditionalnode$139;
assign wirenode$129 = conditionalnode$139;

logic [4:0] zeroextendnode$140;
assign eqnode$130 = wirenode$8 == zeroextendnode$140;

logic [31:0] wirenode$141;
always_ff @ (posedge clock) registernode$131 <= wirenode$141;

logic eqnode$142;
logic [31:0] registernode$143;
logic [31:0] conditionalnode$144;
assign conditionalnode$132 = eqnode$142 ? registernode$143 : conditionalnode$144;

assign zeroextendnode$133 = 4'b1010;

logic [4:0] zeroextendnode$145;
assign eqnode$134 = wirenode$13 == zeroextendnode$145;

logic eqnode$146;
logic [31:0] conditionalnode$147;
assign conditionalnode$135 = eqnode$146 ? registernode$143 : conditionalnode$147;

assign zeroextendnode$136 = 3'b111;

logic [4:0] zeroextendnode$148;
assign eqnode$137 = wirenode$25 == zeroextendnode$148;

logic eqnode$149;
assign andnode$138 = eqnode$149 & wirenode$18;

logic andnode$150;
assign conditionalnode$139 = andnode$150 ? wirenode$11 : registernode$119;

assign zeroextendnode$140 = 4'b1011;

logic [31:0] conditionalnode$151;
assign wirenode$141 = conditionalnode$151;

logic [4:0] zeroextendnode$152;
assign eqnode$142 = wirenode$8 == zeroextendnode$152;

logic [31:0] wirenode$153;
always_ff @ (posedge clock) registernode$143 <= wirenode$153;

logic eqnode$154;
logic [31:0] registernode$155;
logic [31:0] conditionalnode$156;
assign conditionalnode$144 = eqnode$154 ? registernode$155 : conditionalnode$156;

assign zeroextendnode$145 = 4'b1011;

logic [4:0] zeroextendnode$157;
assign eqnode$146 = wirenode$13 == zeroextendnode$157;

logic eqnode$158;
logic [31:0] conditionalnode$159;
assign conditionalnode$147 = eqnode$158 ? registernode$155 : conditionalnode$159;

assign zeroextendnode$148 = 4'b1000;

logic [4:0] zeroextendnode$160;
assign eqnode$149 = wirenode$25 == zeroextendnode$160;

logic eqnode$161;
assign andnode$150 = eqnode$161 & wirenode$18;

logic andnode$162;
assign conditionalnode$151 = andnode$162 ? wirenode$11 : registernode$131;

assign zeroextendnode$152 = 4'b1100;

logic [31:0] conditionalnode$163;
assign wirenode$153 = conditionalnode$163;

logic [4:0] zeroextendnode$164;
assign eqnode$154 = wirenode$8 == zeroextendnode$164;

logic [31:0] wirenode$165;
always_ff @ (posedge clock) registernode$155 <= wirenode$165;

logic eqnode$166;
logic [31:0] registernode$167;
logic [31:0] conditionalnode$168;
assign conditionalnode$156 = eqnode$166 ? registernode$167 : conditionalnode$168;

assign zeroextendnode$157 = 4'b1100;

logic [4:0] zeroextendnode$169;
assign eqnode$158 = wirenode$13 == zeroextendnode$169;

logic eqnode$170;
logic [31:0] conditionalnode$171;
assign conditionalnode$159 = eqnode$170 ? registernode$167 : conditionalnode$171;

assign zeroextendnode$160 = 4'b1001;

logic [4:0] zeroextendnode$172;
assign eqnode$161 = wirenode$25 == zeroextendnode$172;

logic eqnode$173;
assign andnode$162 = eqnode$173 & wirenode$18;

logic andnode$174;
assign conditionalnode$163 = andnode$174 ? wirenode$11 : registernode$143;

assign zeroextendnode$164 = 4'b1101;

logic [31:0] conditionalnode$175;
assign wirenode$165 = conditionalnode$175;

logic [4:0] zeroextendnode$176;
assign eqnode$166 = wirenode$8 == zeroextendnode$176;

logic [31:0] wirenode$177;
always_ff @ (posedge clock) registernode$167 <= wirenode$177;

logic eqnode$178;
logic [31:0] registernode$179;
logic [31:0] conditionalnode$180;
assign conditionalnode$168 = eqnode$178 ? registernode$179 : conditionalnode$180;

assign zeroextendnode$169 = 4'b1101;

logic [4:0] zeroextendnode$181;
assign eqnode$170 = wirenode$13 == zeroextendnode$181;

logic eqnode$182;
logic [31:0] conditionalnode$183;
assign conditionalnode$171 = eqnode$182 ? registernode$179 : conditionalnode$183;

assign zeroextendnode$172 = 4'b1010;

logic [4:0] zeroextendnode$184;
assign eqnode$173 = wirenode$25 == zeroextendnode$184;

logic eqnode$185;
assign andnode$174 = eqnode$185 & wirenode$18;

logic andnode$186;
assign conditionalnode$175 = andnode$186 ? wirenode$11 : registernode$155;

assign zeroextendnode$176 = 4'b1110;

logic [31:0] conditionalnode$187;
assign wirenode$177 = conditionalnode$187;

logic [4:0] zeroextendnode$188;
assign eqnode$178 = wirenode$8 == zeroextendnode$188;

logic [31:0] wirenode$189;
always_ff @ (posedge clock) registernode$179 <= wirenode$189;

logic eqnode$190;
logic [31:0] registernode$191;
logic [31:0] conditionalnode$192;
assign conditionalnode$180 = eqnode$190 ? registernode$191 : conditionalnode$192;

assign zeroextendnode$181 = 4'b1110;

logic [4:0] zeroextendnode$193;
assign eqnode$182 = wirenode$13 == zeroextendnode$193;

logic eqnode$194;
logic [31:0] conditionalnode$195;
assign conditionalnode$183 = eqnode$194 ? registernode$191 : conditionalnode$195;

assign zeroextendnode$184 = 4'b1011;

logic [4:0] zeroextendnode$196;
assign eqnode$185 = wirenode$25 == zeroextendnode$196;

logic eqnode$197;
assign andnode$186 = eqnode$197 & wirenode$18;

logic andnode$198;
assign conditionalnode$187 = andnode$198 ? wirenode$11 : registernode$167;

assign zeroextendnode$188 = 4'b1111;

logic [31:0] conditionalnode$199;
assign wirenode$189 = conditionalnode$199;

assign eqnode$190 = wirenode$8 == 5'b10000;

logic [31:0] wirenode$200;
always_ff @ (posedge clock) registernode$191 <= wirenode$200;

logic eqnode$201;
logic [31:0] registernode$202;
logic [31:0] conditionalnode$203;
assign conditionalnode$192 = eqnode$201 ? registernode$202 : conditionalnode$203;

assign zeroextendnode$193 = 4'b1111;

assign eqnode$194 = wirenode$13 == 5'b10000;

logic eqnode$204;
logic [31:0] conditionalnode$205;
assign conditionalnode$195 = eqnode$204 ? registernode$202 : conditionalnode$205;

assign zeroextendnode$196 = 4'b1100;

logic [4:0] zeroextendnode$206;
assign eqnode$197 = wirenode$25 == zeroextendnode$206;

logic eqnode$207;
assign andnode$198 = eqnode$207 & wirenode$18;

logic andnode$208;
assign conditionalnode$199 = andnode$208 ? wirenode$11 : registernode$179;

logic [31:0] conditionalnode$209;
assign wirenode$200 = conditionalnode$209;

assign eqnode$201 = wirenode$8 == 5'b10001;

logic [31:0] wirenode$210;
always_ff @ (posedge clock) registernode$202 <= wirenode$210;

logic eqnode$211;
logic [31:0] registernode$212;
logic [31:0] conditionalnode$213;
assign conditionalnode$203 = eqnode$211 ? registernode$212 : conditionalnode$213;

assign eqnode$204 = wirenode$13 == 5'b10001;

logic eqnode$214;
logic [31:0] conditionalnode$215;
assign conditionalnode$205 = eqnode$214 ? registernode$212 : conditionalnode$215;

assign zeroextendnode$206 = 4'b1101;

logic [4:0] zeroextendnode$216;
assign eqnode$207 = wirenode$25 == zeroextendnode$216;

logic eqnode$217;
assign andnode$208 = eqnode$217 & wirenode$18;

logic andnode$218;
assign conditionalnode$209 = andnode$218 ? wirenode$11 : registernode$191;

logic [31:0] conditionalnode$219;
assign wirenode$210 = conditionalnode$219;

assign eqnode$211 = wirenode$8 == 5'b10010;

logic [31:0] wirenode$220;
always_ff @ (posedge clock) registernode$212 <= wirenode$220;

logic eqnode$221;
logic [31:0] registernode$222;
logic [31:0] conditionalnode$223;
assign conditionalnode$213 = eqnode$221 ? registernode$222 : conditionalnode$223;

assign eqnode$214 = wirenode$13 == 5'b10010;

logic eqnode$224;
logic [31:0] conditionalnode$225;
assign conditionalnode$215 = eqnode$224 ? registernode$222 : conditionalnode$225;

assign zeroextendnode$216 = 4'b1110;

logic [4:0] zeroextendnode$226;
assign eqnode$217 = wirenode$25 == zeroextendnode$226;

logic eqnode$227;
assign andnode$218 = eqnode$227 & wirenode$18;

logic andnode$228;
assign conditionalnode$219 = andnode$228 ? wirenode$11 : registernode$202;

logic [31:0] conditionalnode$229;
assign wirenode$220 = conditionalnode$229;

assign eqnode$221 = wirenode$8 == 5'b10011;

logic [31:0] wirenode$230;
always_ff @ (posedge clock) registernode$222 <= wirenode$230;

logic eqnode$231;
logic [31:0] registernode$232;
logic [31:0] conditionalnode$233;
assign conditionalnode$223 = eqnode$231 ? registernode$232 : conditionalnode$233;

assign eqnode$224 = wirenode$13 == 5'b10011;

logic eqnode$234;
logic [31:0] conditionalnode$235;
assign conditionalnode$225 = eqnode$234 ? registernode$232 : conditionalnode$235;

assign zeroextendnode$226 = 4'b1111;

assign eqnode$227 = wirenode$25 == 5'b10000;

logic eqnode$236;
assign andnode$228 = eqnode$236 & wirenode$18;

logic andnode$237;
assign conditionalnode$229 = andnode$237 ? wirenode$11 : registernode$212;

logic [31:0] conditionalnode$238;
assign wirenode$230 = conditionalnode$238;

assign eqnode$231 = wirenode$8 == 5'b10100;

logic [31:0] wirenode$239;
always_ff @ (posedge clock) registernode$232 <= wirenode$239;

logic eqnode$240;
logic [31:0] registernode$241;
logic [31:0] conditionalnode$242;
assign conditionalnode$233 = eqnode$240 ? registernode$241 : conditionalnode$242;

assign eqnode$234 = wirenode$13 == 5'b10100;

logic eqnode$243;
logic [31:0] conditionalnode$244;
assign conditionalnode$235 = eqnode$243 ? registernode$241 : conditionalnode$244;

assign eqnode$236 = wirenode$25 == 5'b10001;

logic eqnode$245;
assign andnode$237 = eqnode$245 & wirenode$18;

logic andnode$246;
assign conditionalnode$238 = andnode$246 ? wirenode$11 : registernode$222;

logic [31:0] conditionalnode$247;
assign wirenode$239 = conditionalnode$247;

assign eqnode$240 = wirenode$8 == 5'b10101;

logic [31:0] wirenode$248;
always_ff @ (posedge clock) registernode$241 <= wirenode$248;

logic eqnode$249;
logic [31:0] registernode$250;
logic [31:0] conditionalnode$251;
assign conditionalnode$242 = eqnode$249 ? registernode$250 : conditionalnode$251;

assign eqnode$243 = wirenode$13 == 5'b10101;

logic eqnode$252;
logic [31:0] conditionalnode$253;
assign conditionalnode$244 = eqnode$252 ? registernode$250 : conditionalnode$253;

assign eqnode$245 = wirenode$25 == 5'b10010;

logic eqnode$254;
assign andnode$246 = eqnode$254 & wirenode$18;

logic andnode$255;
assign conditionalnode$247 = andnode$255 ? wirenode$11 : registernode$232;

logic [31:0] conditionalnode$256;
assign wirenode$248 = conditionalnode$256;

assign eqnode$249 = wirenode$8 == 5'b10110;

logic [31:0] wirenode$257;
always_ff @ (posedge clock) registernode$250 <= wirenode$257;

logic eqnode$258;
logic [31:0] registernode$259;
logic [31:0] conditionalnode$260;
assign conditionalnode$251 = eqnode$258 ? registernode$259 : conditionalnode$260;

assign eqnode$252 = wirenode$13 == 5'b10110;

logic eqnode$261;
logic [31:0] conditionalnode$262;
assign conditionalnode$253 = eqnode$261 ? registernode$259 : conditionalnode$262;

assign eqnode$254 = wirenode$25 == 5'b10011;

logic eqnode$263;
assign andnode$255 = eqnode$263 & wirenode$18;

logic andnode$264;
assign conditionalnode$256 = andnode$264 ? wirenode$11 : registernode$241;

logic [31:0] conditionalnode$265;
assign wirenode$257 = conditionalnode$265;

assign eqnode$258 = wirenode$8 == 5'b10111;

logic [31:0] wirenode$266;
always_ff @ (posedge clock) registernode$259 <= wirenode$266;

logic eqnode$267;
logic [31:0] registernode$268;
logic [31:0] conditionalnode$269;
assign conditionalnode$260 = eqnode$267 ? registernode$268 : conditionalnode$269;

assign eqnode$261 = wirenode$13 == 5'b10111;

logic eqnode$270;
logic [31:0] conditionalnode$271;
assign conditionalnode$262 = eqnode$270 ? registernode$268 : conditionalnode$271;

assign eqnode$263 = wirenode$25 == 5'b10100;

logic eqnode$272;
assign andnode$264 = eqnode$272 & wirenode$18;

logic andnode$273;
assign conditionalnode$265 = andnode$273 ? wirenode$11 : registernode$250;

logic [31:0] conditionalnode$274;
assign wirenode$266 = conditionalnode$274;

assign eqnode$267 = wirenode$8 == 5'b11000;

logic [31:0] wirenode$275;
always_ff @ (posedge clock) registernode$268 <= wirenode$275;

logic eqnode$276;
logic [31:0] registernode$277;
logic [31:0] conditionalnode$278;
assign conditionalnode$269 = eqnode$276 ? registernode$277 : conditionalnode$278;

assign eqnode$270 = wirenode$13 == 5'b11000;

logic eqnode$279;
logic [31:0] conditionalnode$280;
assign conditionalnode$271 = eqnode$279 ? registernode$277 : conditionalnode$280;

assign eqnode$272 = wirenode$25 == 5'b10101;

logic eqnode$281;
assign andnode$273 = eqnode$281 & wirenode$18;

logic andnode$282;
assign conditionalnode$274 = andnode$282 ? wirenode$11 : registernode$259;

logic [31:0] conditionalnode$283;
assign wirenode$275 = conditionalnode$283;

assign eqnode$276 = wirenode$8 == 5'b11001;

logic [31:0] wirenode$284;
always_ff @ (posedge clock) registernode$277 <= wirenode$284;

logic eqnode$285;
logic [31:0] registernode$286;
logic [31:0] conditionalnode$287;
assign conditionalnode$278 = eqnode$285 ? registernode$286 : conditionalnode$287;

assign eqnode$279 = wirenode$13 == 5'b11001;

logic eqnode$288;
logic [31:0] conditionalnode$289;
assign conditionalnode$280 = eqnode$288 ? registernode$286 : conditionalnode$289;

assign eqnode$281 = wirenode$25 == 5'b10110;

logic eqnode$290;
assign andnode$282 = eqnode$290 & wirenode$18;

logic andnode$291;
assign conditionalnode$283 = andnode$291 ? wirenode$11 : registernode$268;

logic [31:0] conditionalnode$292;
assign wirenode$284 = conditionalnode$292;

assign eqnode$285 = wirenode$8 == 5'b11010;

logic [31:0] wirenode$293;
always_ff @ (posedge clock) registernode$286 <= wirenode$293;

logic eqnode$294;
logic [31:0] registernode$295;
logic [31:0] conditionalnode$296;
assign conditionalnode$287 = eqnode$294 ? registernode$295 : conditionalnode$296;

assign eqnode$288 = wirenode$13 == 5'b11010;

logic eqnode$297;
logic [31:0] conditionalnode$298;
assign conditionalnode$289 = eqnode$297 ? registernode$295 : conditionalnode$298;

assign eqnode$290 = wirenode$25 == 5'b10111;

logic eqnode$299;
assign andnode$291 = eqnode$299 & wirenode$18;

logic andnode$300;
assign conditionalnode$292 = andnode$300 ? wirenode$11 : registernode$277;

logic [31:0] conditionalnode$301;
assign wirenode$293 = conditionalnode$301;

assign eqnode$294 = wirenode$8 == 5'b11011;

logic [31:0] wirenode$302;
always_ff @ (posedge clock) registernode$295 <= wirenode$302;

logic eqnode$303;
logic [31:0] registernode$304;
logic [31:0] conditionalnode$305;
assign conditionalnode$296 = eqnode$303 ? registernode$304 : conditionalnode$305;

assign eqnode$297 = wirenode$13 == 5'b11011;

logic eqnode$306;
logic [31:0] conditionalnode$307;
assign conditionalnode$298 = eqnode$306 ? registernode$304 : conditionalnode$307;

assign eqnode$299 = wirenode$25 == 5'b11000;

logic eqnode$308;
assign andnode$300 = eqnode$308 & wirenode$18;

logic andnode$309;
assign conditionalnode$301 = andnode$309 ? wirenode$11 : registernode$286;

logic [31:0] conditionalnode$310;
assign wirenode$302 = conditionalnode$310;

assign eqnode$303 = wirenode$8 == 5'b11100;

logic [31:0] wirenode$311;
always_ff @ (posedge clock) registernode$304 <= wirenode$311;

logic eqnode$312;
logic [31:0] registernode$313;
logic [31:0] conditionalnode$314;
assign conditionalnode$305 = eqnode$312 ? registernode$313 : conditionalnode$314;

assign eqnode$306 = wirenode$13 == 5'b11100;

logic eqnode$315;
logic [31:0] conditionalnode$316;
assign conditionalnode$307 = eqnode$315 ? registernode$313 : conditionalnode$316;

assign eqnode$308 = wirenode$25 == 5'b11001;

logic eqnode$317;
assign andnode$309 = eqnode$317 & wirenode$18;

logic andnode$318;
assign conditionalnode$310 = andnode$318 ? wirenode$11 : registernode$295;

logic [31:0] conditionalnode$319;
assign wirenode$311 = conditionalnode$319;

assign eqnode$312 = wirenode$8 == 5'b11101;

logic [31:0] wirenode$320;
always_ff @ (posedge clock) registernode$313 <= wirenode$320;

logic eqnode$321;
logic [31:0] registernode$322;
logic [31:0] conditionalnode$323;
assign conditionalnode$314 = eqnode$321 ? registernode$322 : conditionalnode$323;

assign eqnode$315 = wirenode$13 == 5'b11101;

logic eqnode$324;
logic [31:0] conditionalnode$325;
assign conditionalnode$316 = eqnode$324 ? registernode$322 : conditionalnode$325;

assign eqnode$317 = wirenode$25 == 5'b11010;

logic eqnode$326;
assign andnode$318 = eqnode$326 & wirenode$18;

logic andnode$327;
assign conditionalnode$319 = andnode$327 ? wirenode$11 : registernode$304;

logic [31:0] conditionalnode$328;
assign wirenode$320 = conditionalnode$328;

assign eqnode$321 = wirenode$8 == 5'b11110;

logic [31:0] wirenode$329;
always_ff @ (posedge clock) registernode$322 <= wirenode$329;

logic eqnode$330;
logic [31:0] registernode$331;
logic [31:0] repeatnode$332;
assign conditionalnode$323 = eqnode$330 ? registernode$331 : repeatnode$332;

assign eqnode$324 = wirenode$13 == 5'b11110;

logic eqnode$333;
logic [31:0] repeatnode$334;
assign conditionalnode$325 = eqnode$333 ? registernode$331 : repeatnode$334;

assign eqnode$326 = wirenode$25 == 5'b11011;

logic eqnode$335;
assign andnode$327 = eqnode$335 & wirenode$18;

logic andnode$336;
assign conditionalnode$328 = andnode$336 ? wirenode$11 : registernode$313;

logic [31:0] conditionalnode$337;
assign wirenode$329 = conditionalnode$337;

assign eqnode$330 = wirenode$8 == 5'b11111;

logic [31:0] wirenode$338;
always_ff @ (posedge clock) registernode$331 <= wirenode$338;

assign repeatnode$332 = {32{1'bX}};

assign eqnode$333 = wirenode$13 == 5'b11111;

assign repeatnode$334 = {32{1'bX}};

assign eqnode$335 = wirenode$25 == 5'b11100;

logic eqnode$339;
assign andnode$336 = eqnode$339 & wirenode$18;

logic andnode$340;
assign conditionalnode$337 = andnode$340 ? wirenode$11 : registernode$322;

logic [31:0] conditionalnode$341;
assign wirenode$338 = conditionalnode$341;

assign eqnode$339 = wirenode$25 == 5'b11101;

logic eqnode$342;
assign andnode$340 = eqnode$342 & wirenode$18;

logic andnode$343;
assign conditionalnode$341 = andnode$343 ? wirenode$11 : registernode$331;

assign eqnode$342 = wirenode$25 == 5'b11110;

logic eqnode$344;
assign andnode$343 = eqnode$344 & wirenode$18;

assign eqnode$344 = wirenode$25 == 5'b11111;

endmodule
